module USFFT64_2B_RING(CLK, CLK_C, RST, RST_C, ED, ED_C, START, START_C, SHIFT, SHIFT_C, DR, DR_C, DI, DI_C, RDY, RDY_C, OVF1, OVF1_C, OVF2, OVF2_C,
     ADDR, ADDR_C, DOR, DOR_C, DOI, DOI_C, dft_shift_enable, dft_shift_enable_C, dft_scan_input_1, dft_scan_input_1_C,
     dft_scan_input_2, dft_scan_input_2_C, dft_scan_output_1, dft_scan_output_1_C, dft_scan_output_2, dft_scan_output_2_C);
  
  input CLK, RST, ED, START, dft_shift_enable, dft_scan_input_1, dft_scan_input_2;
  input [3:0] SHIFT;
  input [15:0] DR, DI;
  output RDY, OVF1, OVF2, dft_scan_output_1, dft_scan_output_2;
  output [5:0] ADDR;
  output [18:0] DOR, DOI;

  output CLK_C, RST_C, ED_C, START_C, dft_shift_enable_C, dft_scan_input_1_C, dft_scan_input_2_C;
  output [3:0] SHIFT_C;
  output [15:0] DR_C, DI_C;
  input RDY_C, OVF1_C, OVF2_C, dft_scan_output_1_C, dft_scan_output_2_C;
  input [5:0] ADDR_C;
  input [18:0] DOR_C, DOI_C;

  wire VDD, VDDO, VDDR, GNDR, GNDO;

  ICF PAD_CLK     (.PAD(CLK),       .Y(CLK_C),      .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_RST     (.PAD(RST),       .Y(RST_C),      .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_ED      (.PAD(ED),        .Y(ED_C),       .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_START   (.PAD(START),     .Y(START_C),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_SHIFT_0 (.PAD(SHIFT[0]),  .Y(SHIFT_C[0]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_SHIFT_1 (.PAD(SHIFT[1]),  .Y(SHIFT_C[1]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_SHIFT_2 (.PAD(SHIFT[2]),  .Y(SHIFT_C[2]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_SHIFT_3 (.PAD(SHIFT[3]),  .Y(SHIFT_C[3]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_0    (.PAD(DR[0]),     .Y(DR_C[0]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_1    (.PAD(DR[1]),     .Y(DR_C[1]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_2    (.PAD(DR[2]),     .Y(DR_C[2]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_3    (.PAD(DR[3]),     .Y(DR_C[3]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_4    (.PAD(DR[4]),     .Y(DR_C[4]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_5    (.PAD(DR[5]),     .Y(DR_C[5]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_6    (.PAD(DR[6]),     .Y(DR_C[6]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_7    (.PAD(DR[7]),     .Y(DR_C[7]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_8    (.PAD(DR[8]),     .Y(DR_C[8]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_9    (.PAD(DR[9]),     .Y(DR_C[9]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_10   (.PAD(DR[10]),    .Y(DR_C[10]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_11   (.PAD(DR[11]),    .Y(DR_C[11]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_12   (.PAD(DR[12]),    .Y(DR_C[12]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_13   (.PAD(DR[13]),    .Y(DR_C[13]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_14   (.PAD(DR[14]),    .Y(DR_C[14]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DR_15   (.PAD(DR[15]),    .Y(DR_C[15]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_0    (.PAD(DI[0]),     .Y(DI_C[0]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_1    (.PAD(DI[1]),     .Y(DI_C[1]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_2    (.PAD(DI[2]),     .Y(DI_C[2]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_3    (.PAD(DI[3]),     .Y(DI_C[3]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_4    (.PAD(DI[4]),     .Y(DI_C[4]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_5    (.PAD(DI[5]),     .Y(DI_C[5]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_6    (.PAD(DI[6]),     .Y(DI_C[6]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_7    (.PAD(DI[7]),     .Y(DI_C[7]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_8    (.PAD(DI[8]),     .Y(DI_C[8]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_9    (.PAD(DI[9]),     .Y(DI_C[9]),    .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_10   (.PAD(DI[10]),    .Y(DI_C[10]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_11   (.PAD(DI[11]),    .Y(DI_C[11]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_12   (.PAD(DI[12]),    .Y(DI_C[12]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_13   (.PAD(DI[13]),    .Y(DI_C[13]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_14   (.PAD(DI[14]),    .Y(DI_C[14]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DI_15   (.PAD(DI[15]),    .Y(DI_C[15]),   .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));

  // Outputs
  BT8SF PAD_RDY  (.A(RDY_C),  .EN(1'b0), .PAD(RDY),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_OVF1 (.A(OVF1_C), .EN(1'b0), .PAD(OVF1), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_OVF2 (.A(OVF2_C), .EN(1'b0), .PAD(OVF2), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DFT_SCAN_OUTPUT_1 (.A(dft_scan_output_1_C), .EN(1'b0), .PAD(dft_scan_output_1), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DFT_SCAN_OUTPUT_2 (.A(dft_scan_output_2_C), .EN(1'b0), .PAD(dft_scan_output_2), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));

  // Inputs
  ICF PAD_DFT_SHIFT_ENABLE (.PAD(dft_shift_enable), .Y(dft_shift_enable_C), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DFT_SCAN_INPUT_1 (.PAD(dft_scan_input_1), .Y(dft_scan_input_1_C), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  ICF PAD_DFT_SCAN_INPUT_2 (.PAD(dft_scan_input_2), .Y(dft_scan_input_2_C), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));

  // ADDR (output)
  BT8SF PAD_ADDR_0 (.A(ADDR_C[0]), .EN(1'b0),.PAD(ADDR[0]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_ADDR_1 (.A(ADDR_C[1]), .EN(1'b0),.PAD(ADDR[1]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_ADDR_2 (.A(ADDR_C[2]), .EN(1'b0),.PAD(ADDR[2]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_ADDR_3 (.A(ADDR_C[3]), .EN(1'b0),.PAD(ADDR[3]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_ADDR_4 (.A(ADDR_C[4]), .EN(1'b0),.PAD(ADDR[4]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_ADDR_5 (.A(ADDR_C[5]), .EN(1'b0),.PAD(ADDR[5]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));

  // DOR (output)
  BT8SF PAD_DOR_0  (.A(DOR_C[0]),  .EN(1'b0),.PAD(DOR[0]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_1  (.A(DOR_C[1]),  .EN(1'b0),.PAD(DOR[1]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_2  (.A(DOR_C[2]),  .EN(1'b0),.PAD(DOR[2]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_3  (.A(DOR_C[3]),  .EN(1'b0),.PAD(DOR[3]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_4  (.A(DOR_C[4]),  .EN(1'b0),.PAD(DOR[4]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_5  (.A(DOR_C[5]),  .EN(1'b0),.PAD(DOR[5]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_6  (.A(DOR_C[6]),  .EN(1'b0),.PAD(DOR[6]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_7  (.A(DOR_C[7]),  .EN(1'b0),.PAD(DOR[7]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_8  (.A(DOR_C[8]),  .EN(1'b0),.PAD(DOR[8]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_9  (.A(DOR_C[9]),  .EN(1'b0),.PAD(DOR[9]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_10 (.A(DOR_C[10]), .EN(1'b0),.PAD(DOR[10]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_11 (.A(DOR_C[11]), .EN(1'b0),.PAD(DOR[11]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_12 (.A(DOR_C[12]), .EN(1'b0),.PAD(DOR[12]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_13 (.A(DOR_C[13]), .EN(1'b0),.PAD(DOR[13]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_14 (.A(DOR_C[14]), .EN(1'b0),.PAD(DOR[14]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_15 (.A(DOR_C[15]), .EN(1'b0),.PAD(DOR[15]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_16 (.A(DOR_C[16]), .EN(1'b0),.PAD(DOR[16]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_17 (.A(DOR_C[17]), .EN(1'b0),.PAD(DOR[17]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOR_18 (.A(DOR_C[18]), .EN(1'b0),.PAD(DOR[18]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));

  // DOI (output)
  BT8SF PAD_DOI_0  (.A(DOI_C[0]),  .EN(1'b0),.PAD(DOI[0]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_1  (.A(DOI_C[1]),  .EN(1'b0),.PAD(DOI[1]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_2  (.A(DOI_C[2]),  .EN(1'b0),.PAD(DOI[2]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_3  (.A(DOI_C[3]),  .EN(1'b0),.PAD(DOI[3]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_4  (.A(DOI_C[4]),  .EN(1'b0),.PAD(DOI[4]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_5  (.A(DOI_C[5]),  .EN(1'b0),.PAD(DOI[5]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_6  (.A(DOI_C[6]),  .EN(1'b0),.PAD(DOI[6]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_7  (.A(DOI_C[7]),  .EN(1'b0),.PAD(DOI[7]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_8  (.A(DOI_C[8]),  .EN(1'b0),.PAD(DOI[8]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_9  (.A(DOI_C[9]),  .EN(1'b0),.PAD(DOI[9]),  .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_10 (.A(DOI_C[10]), .EN(1'b0),.PAD(DOI[10]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_11 (.A(DOI_C[11]), .EN(1'b0),.PAD(DOI[11]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_12 (.A(DOI_C[12]), .EN(1'b0),.PAD(DOI[12]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_13 (.A(DOI_C[13]), .EN(1'b0),.PAD(DOI[13]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_14 (.A(DOI_C[14]), .EN(1'b0),.PAD(DOI[14]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_15 (.A(DOI_C[15]), .EN(1'b0),.PAD(DOI[15]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_16 (.A(DOI_C[16]), .EN(1'b0),.PAD(DOI[16]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_17 (.A(DOI_C[17]), .EN(1'b0),.PAD(DOI[17]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));
  BT8SF PAD_DOI_18 (.A(DOI_C[18]), .EN(1'b0),.PAD(DOI[18]), .VDD(VDD), .VDDO(VDDO), .VDDR(VDDR), .GNDR(GNDR), .GNDO(GNDO));

  CORNERF CORNER_TL (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
  CORNERF CORNER_TR (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
  CORNERF CORNER_BL (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
  CORNERF CORNER_BR (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));

  VDDIPADF VDD_C_N (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
  VDDIPADF VDD_C_S (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
  VDDIPADF VDD_C_W (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR)); 
  VDDIPADF VDD_C_E (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
  GNDIPADF GND_C_N (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
  GNDIPADF GND_C_S (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
  GNDIPADF GND_C_W (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
  GNDIPADF GND_C_E (.GNDO(GNDO),.GNDR(GNDR),.VDD(VDD),.VDDO(VDDO),.VDDR(VDDR));
    
  
 endmodule

